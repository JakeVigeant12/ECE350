module(data,inverted_data);
input [31:0] data;
output [31:0] inverted_data;
not not0(inverted_data[0], data[0]);
not not1(inverted_data[1], data[1]);
not not2(inverted_data[2], data[2]);
not not3(inverted_data[3], data[3]);
not not4(inverted_data[4], data[4]);
not not5(inverted_data[5], data[5]);
not not6(inverted_data[6], data[6]);
not not7(inverted_data[7], data[7]);
not not8(inverted_data[8], data[8]);
not not9(inverted_data[9], data[9]);
not not10(inverted_data[10], data[10]);
not not11(inverted_data[11], data[11]);
not not12(inverted_data[12], data[12]);
not not13(inverted_data[13], data[13]);
not not14(inverted_data[14], data[14]);
not not15(inverted_data[15], data[15]);
not not16(inverted_data[16], data[16]);
not not17(inverted_data[17], data[17]);
not not18(inverted_data[18], data[18]);
not not19(inverted_data[19], data[19]);
not not20(inverted_data[20], data[20]);
not not21(inverted_data[21], data[21]);
not not22(inverted_data[22], data[22]);
not not23(inverted_data[23], data[23]);
not not24(inverted_data[24], data[24]);
not not25(inverted_data[25], data[25]);
not not26(inverted_data[26], data[26]);
not not27(inverted_data[27], data[27]);
not not28(inverted_data[28], data[28]);
not not29(inverted_data[29], data[29]);
not not30(inverted_data[30], data[30]);
not not31(inverted_data[31], data[31]);
endmodule